module RF( // @[:RF.fir@3.2]
  input        clock, // @[:RF.fir@4.4]
  input        reset, // @[:RF.fir@5.4]
  input        io_control_internal_wEnable_0, // @[:RF.fir@6.4]
  input        io_control_internal_rEnable_0, // @[:RF.fir@6.4]
  input  [4:0] io_control_internal_wAddr_0, // @[:RF.fir@6.4]
  input  [4:0] io_control_internal_rAddr_0, // @[:RF.fir@6.4]
  input        io_control_internal_bpSel_0_0, // @[:RF.fir@6.4]
  input        io_control_external_wEnable_0, // @[:RF.fir@6.4]
  input        io_control_external_rEnable_0, // @[:RF.fir@6.4]
  input  [4:0] io_control_external_wAddr_0, // @[:RF.fir@6.4]
  input  [4:0] io_control_external_rAddr_0, // @[:RF.fir@6.4]
  input        io_control_external_bpSel_0_0, // @[:RF.fir@6.4]
  input  [7:0] io_wInternal_0, // @[:RF.fir@6.4]
  input  [7:0] io_wExternal_0, // @[:RF.fir@6.4]
  output [7:0] io_rInternal_0, // @[:RF.fir@6.4]
  output [7:0] io_rExternal_0 // @[:RF.fir@6.4]
);
  reg [7:0] dataRegister_0; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_0;
  reg [7:0] dataRegister_1; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_1;
  reg [7:0] dataRegister_2; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_2;
  reg [7:0] dataRegister_3; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_3;
  reg [7:0] dataRegister_4; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_4;
  reg [7:0] dataRegister_5; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_5;
  reg [7:0] dataRegister_6; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_6;
  reg [7:0] dataRegister_7; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_7;
  reg [7:0] dataRegister_8; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_8;
  reg [7:0] dataRegister_9; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_9;
  reg [7:0] dataRegister_10; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_10;
  reg [7:0] dataRegister_11; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_11;
  reg [7:0] dataRegister_12; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_12;
  reg [7:0] dataRegister_13; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_13;
  reg [7:0] dataRegister_14; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_14;
  reg [7:0] dataRegister_15; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_15;
  reg [7:0] dataRegister_16; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_16;
  reg [7:0] dataRegister_17; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_17;
  reg [7:0] dataRegister_18; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_18;
  reg [7:0] dataRegister_19; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_19;
  reg [7:0] dataRegister_20; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_20;
  reg [7:0] dataRegister_21; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_21;
  reg [7:0] dataRegister_22; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_22;
  reg [7:0] dataRegister_23; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_23;
  reg [7:0] dataRegister_24; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_24;
  reg [7:0] dataRegister_25; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_25;
  reg [7:0] dataRegister_26; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_26;
  reg [7:0] dataRegister_27; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_27;
  reg [7:0] dataRegister_28; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_28;
  reg [7:0] dataRegister_29; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_29;
  reg [7:0] dataRegister_30; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_30;
  reg [7:0] dataRegister_31; // @[PE.scala 76:21:RF.fir@41.4]
  reg [31:0] _RAND_31;
  reg [7:0] bpRegisterInt_0; // @[PE.scala 81:21:RF.fir@44.4]
  reg [31:0] _RAND_32;
  reg [7:0] bpRegisterExt_0; // @[PE.scala 83:21:RF.fir@47.4]
  reg [31:0] _RAND_33;
  wire [7:0] _GEN_131; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_132; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_133; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_134; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_135; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_136; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_137; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_138; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_139; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_140; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_141; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_142; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_143; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_144; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_145; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_146; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_147; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_148; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_149; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_150; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_151; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_152; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_153; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_154; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_155; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_156; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_157; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_158; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_159; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_160; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_161; // @[PE.scala 108:37:RF.fir@63.8]
  wire [7:0] _GEN_162; // @[PE.scala 104:78:RF.fir@59.6]
  wire [7:0] _GEN_165; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_166; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_167; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_168; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_169; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_170; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_171; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_172; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_173; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_174; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_175; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_176; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_177; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_178; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_179; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_180; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_181; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_182; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_183; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_184; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_185; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_186; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_187; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_188; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_189; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_190; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_191; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_192; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_193; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_194; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_195; // @[PE.scala 127:37:RF.fir@76.8]
  wire [7:0] _GEN_196; // @[PE.scala 123:78:RF.fir@72.6]
  assign _GEN_131 = 5'h1 == io_control_internal_rAddr_0 ? $signed(dataRegister_1) : $signed(dataRegister_0); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_132 = 5'h2 == io_control_internal_rAddr_0 ? $signed(dataRegister_2) : $signed(_GEN_131); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_133 = 5'h3 == io_control_internal_rAddr_0 ? $signed(dataRegister_3) : $signed(_GEN_132); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_134 = 5'h4 == io_control_internal_rAddr_0 ? $signed(dataRegister_4) : $signed(_GEN_133); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_135 = 5'h5 == io_control_internal_rAddr_0 ? $signed(dataRegister_5) : $signed(_GEN_134); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_136 = 5'h6 == io_control_internal_rAddr_0 ? $signed(dataRegister_6) : $signed(_GEN_135); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_137 = 5'h7 == io_control_internal_rAddr_0 ? $signed(dataRegister_7) : $signed(_GEN_136); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_138 = 5'h8 == io_control_internal_rAddr_0 ? $signed(dataRegister_8) : $signed(_GEN_137); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_139 = 5'h9 == io_control_internal_rAddr_0 ? $signed(dataRegister_9) : $signed(_GEN_138); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_140 = 5'ha == io_control_internal_rAddr_0 ? $signed(dataRegister_10) : $signed(_GEN_139); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_141 = 5'hb == io_control_internal_rAddr_0 ? $signed(dataRegister_11) : $signed(_GEN_140); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_142 = 5'hc == io_control_internal_rAddr_0 ? $signed(dataRegister_12) : $signed(_GEN_141); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_143 = 5'hd == io_control_internal_rAddr_0 ? $signed(dataRegister_13) : $signed(_GEN_142); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_144 = 5'he == io_control_internal_rAddr_0 ? $signed(dataRegister_14) : $signed(_GEN_143); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_145 = 5'hf == io_control_internal_rAddr_0 ? $signed(dataRegister_15) : $signed(_GEN_144); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_146 = 5'h10 == io_control_internal_rAddr_0 ? $signed(dataRegister_16) : $signed(_GEN_145); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_147 = 5'h11 == io_control_internal_rAddr_0 ? $signed(dataRegister_17) : $signed(_GEN_146); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_148 = 5'h12 == io_control_internal_rAddr_0 ? $signed(dataRegister_18) : $signed(_GEN_147); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_149 = 5'h13 == io_control_internal_rAddr_0 ? $signed(dataRegister_19) : $signed(_GEN_148); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_150 = 5'h14 == io_control_internal_rAddr_0 ? $signed(dataRegister_20) : $signed(_GEN_149); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_151 = 5'h15 == io_control_internal_rAddr_0 ? $signed(dataRegister_21) : $signed(_GEN_150); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_152 = 5'h16 == io_control_internal_rAddr_0 ? $signed(dataRegister_22) : $signed(_GEN_151); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_153 = 5'h17 == io_control_internal_rAddr_0 ? $signed(dataRegister_23) : $signed(_GEN_152); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_154 = 5'h18 == io_control_internal_rAddr_0 ? $signed(dataRegister_24) : $signed(_GEN_153); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_155 = 5'h19 == io_control_internal_rAddr_0 ? $signed(dataRegister_25) : $signed(_GEN_154); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_156 = 5'h1a == io_control_internal_rAddr_0 ? $signed(dataRegister_26) : $signed(_GEN_155); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_157 = 5'h1b == io_control_internal_rAddr_0 ? $signed(dataRegister_27) : $signed(_GEN_156); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_158 = 5'h1c == io_control_internal_rAddr_0 ? $signed(dataRegister_28) : $signed(_GEN_157); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_159 = 5'h1d == io_control_internal_rAddr_0 ? $signed(dataRegister_29) : $signed(_GEN_158); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_160 = 5'h1e == io_control_internal_rAddr_0 ? $signed(dataRegister_30) : $signed(_GEN_159); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_161 = 5'h1f == io_control_internal_rAddr_0 ? $signed(dataRegister_31) : $signed(_GEN_160); // @[PE.scala 108:37:RF.fir@63.8]
  assign _GEN_162 = io_control_internal_bpSel_0_0 ? $signed(bpRegisterExt_0) : $signed(_GEN_161); // @[PE.scala 104:78:RF.fir@59.6]
  assign _GEN_165 = 5'h1 == io_control_external_rAddr_0 ? $signed(dataRegister_1) : $signed(dataRegister_0); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_166 = 5'h2 == io_control_external_rAddr_0 ? $signed(dataRegister_2) : $signed(_GEN_165); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_167 = 5'h3 == io_control_external_rAddr_0 ? $signed(dataRegister_3) : $signed(_GEN_166); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_168 = 5'h4 == io_control_external_rAddr_0 ? $signed(dataRegister_4) : $signed(_GEN_167); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_169 = 5'h5 == io_control_external_rAddr_0 ? $signed(dataRegister_5) : $signed(_GEN_168); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_170 = 5'h6 == io_control_external_rAddr_0 ? $signed(dataRegister_6) : $signed(_GEN_169); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_171 = 5'h7 == io_control_external_rAddr_0 ? $signed(dataRegister_7) : $signed(_GEN_170); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_172 = 5'h8 == io_control_external_rAddr_0 ? $signed(dataRegister_8) : $signed(_GEN_171); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_173 = 5'h9 == io_control_external_rAddr_0 ? $signed(dataRegister_9) : $signed(_GEN_172); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_174 = 5'ha == io_control_external_rAddr_0 ? $signed(dataRegister_10) : $signed(_GEN_173); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_175 = 5'hb == io_control_external_rAddr_0 ? $signed(dataRegister_11) : $signed(_GEN_174); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_176 = 5'hc == io_control_external_rAddr_0 ? $signed(dataRegister_12) : $signed(_GEN_175); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_177 = 5'hd == io_control_external_rAddr_0 ? $signed(dataRegister_13) : $signed(_GEN_176); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_178 = 5'he == io_control_external_rAddr_0 ? $signed(dataRegister_14) : $signed(_GEN_177); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_179 = 5'hf == io_control_external_rAddr_0 ? $signed(dataRegister_15) : $signed(_GEN_178); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_180 = 5'h10 == io_control_external_rAddr_0 ? $signed(dataRegister_16) : $signed(_GEN_179); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_181 = 5'h11 == io_control_external_rAddr_0 ? $signed(dataRegister_17) : $signed(_GEN_180); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_182 = 5'h12 == io_control_external_rAddr_0 ? $signed(dataRegister_18) : $signed(_GEN_181); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_183 = 5'h13 == io_control_external_rAddr_0 ? $signed(dataRegister_19) : $signed(_GEN_182); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_184 = 5'h14 == io_control_external_rAddr_0 ? $signed(dataRegister_20) : $signed(_GEN_183); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_185 = 5'h15 == io_control_external_rAddr_0 ? $signed(dataRegister_21) : $signed(_GEN_184); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_186 = 5'h16 == io_control_external_rAddr_0 ? $signed(dataRegister_22) : $signed(_GEN_185); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_187 = 5'h17 == io_control_external_rAddr_0 ? $signed(dataRegister_23) : $signed(_GEN_186); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_188 = 5'h18 == io_control_external_rAddr_0 ? $signed(dataRegister_24) : $signed(_GEN_187); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_189 = 5'h19 == io_control_external_rAddr_0 ? $signed(dataRegister_25) : $signed(_GEN_188); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_190 = 5'h1a == io_control_external_rAddr_0 ? $signed(dataRegister_26) : $signed(_GEN_189); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_191 = 5'h1b == io_control_external_rAddr_0 ? $signed(dataRegister_27) : $signed(_GEN_190); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_192 = 5'h1c == io_control_external_rAddr_0 ? $signed(dataRegister_28) : $signed(_GEN_191); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_193 = 5'h1d == io_control_external_rAddr_0 ? $signed(dataRegister_29) : $signed(_GEN_192); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_194 = 5'h1e == io_control_external_rAddr_0 ? $signed(dataRegister_30) : $signed(_GEN_193); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_195 = 5'h1f == io_control_external_rAddr_0 ? $signed(dataRegister_31) : $signed(_GEN_194); // @[PE.scala 127:37:RF.fir@76.8]
  assign _GEN_196 = io_control_external_bpSel_0_0 ? $signed(bpRegisterInt_0) : $signed(_GEN_195); // @[PE.scala 123:78:RF.fir@72.6]
  assign io_rInternal_0 = io_control_internal_rEnable_0 ? $signed(_GEN_162) : $signed(8'sh0);
  assign io_rExternal_0 = io_control_external_rEnable_0 ? $signed(_GEN_196) : $signed(8'sh0);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  dataRegister_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  dataRegister_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  dataRegister_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  dataRegister_3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  dataRegister_4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  dataRegister_5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  dataRegister_6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  dataRegister_7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  dataRegister_8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  dataRegister_9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  dataRegister_10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  dataRegister_11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  dataRegister_12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  dataRegister_13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  dataRegister_14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  dataRegister_15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  dataRegister_16 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  dataRegister_17 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  dataRegister_18 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  dataRegister_19 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  dataRegister_20 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  dataRegister_21 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  dataRegister_22 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  dataRegister_23 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  dataRegister_24 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  dataRegister_25 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  dataRegister_26 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  dataRegister_27 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  dataRegister_28 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  dataRegister_29 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  dataRegister_30 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  dataRegister_31 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  bpRegisterInt_0 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  bpRegisterExt_0 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      dataRegister_0 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h0 == io_control_external_wAddr_0) begin
          dataRegister_0 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h0 == io_control_internal_wAddr_0) begin
              dataRegister_0 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h0 == io_control_internal_wAddr_0) begin
            dataRegister_0 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_1 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h1 == io_control_external_wAddr_0) begin
          dataRegister_1 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h1 == io_control_internal_wAddr_0) begin
              dataRegister_1 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h1 == io_control_internal_wAddr_0) begin
            dataRegister_1 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_2 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h2 == io_control_external_wAddr_0) begin
          dataRegister_2 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h2 == io_control_internal_wAddr_0) begin
              dataRegister_2 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h2 == io_control_internal_wAddr_0) begin
            dataRegister_2 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_3 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h3 == io_control_external_wAddr_0) begin
          dataRegister_3 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h3 == io_control_internal_wAddr_0) begin
              dataRegister_3 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h3 == io_control_internal_wAddr_0) begin
            dataRegister_3 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_4 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h4 == io_control_external_wAddr_0) begin
          dataRegister_4 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h4 == io_control_internal_wAddr_0) begin
              dataRegister_4 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h4 == io_control_internal_wAddr_0) begin
            dataRegister_4 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_5 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h5 == io_control_external_wAddr_0) begin
          dataRegister_5 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h5 == io_control_internal_wAddr_0) begin
              dataRegister_5 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h5 == io_control_internal_wAddr_0) begin
            dataRegister_5 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_6 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h6 == io_control_external_wAddr_0) begin
          dataRegister_6 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h6 == io_control_internal_wAddr_0) begin
              dataRegister_6 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h6 == io_control_internal_wAddr_0) begin
            dataRegister_6 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_7 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h7 == io_control_external_wAddr_0) begin
          dataRegister_7 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h7 == io_control_internal_wAddr_0) begin
              dataRegister_7 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h7 == io_control_internal_wAddr_0) begin
            dataRegister_7 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_8 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h8 == io_control_external_wAddr_0) begin
          dataRegister_8 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h8 == io_control_internal_wAddr_0) begin
              dataRegister_8 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h8 == io_control_internal_wAddr_0) begin
            dataRegister_8 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_9 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h9 == io_control_external_wAddr_0) begin
          dataRegister_9 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h9 == io_control_internal_wAddr_0) begin
              dataRegister_9 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h9 == io_control_internal_wAddr_0) begin
            dataRegister_9 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_10 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'ha == io_control_external_wAddr_0) begin
          dataRegister_10 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'ha == io_control_internal_wAddr_0) begin
              dataRegister_10 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'ha == io_control_internal_wAddr_0) begin
            dataRegister_10 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_11 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'hb == io_control_external_wAddr_0) begin
          dataRegister_11 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'hb == io_control_internal_wAddr_0) begin
              dataRegister_11 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'hb == io_control_internal_wAddr_0) begin
            dataRegister_11 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_12 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'hc == io_control_external_wAddr_0) begin
          dataRegister_12 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'hc == io_control_internal_wAddr_0) begin
              dataRegister_12 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'hc == io_control_internal_wAddr_0) begin
            dataRegister_12 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_13 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'hd == io_control_external_wAddr_0) begin
          dataRegister_13 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'hd == io_control_internal_wAddr_0) begin
              dataRegister_13 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'hd == io_control_internal_wAddr_0) begin
            dataRegister_13 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_14 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'he == io_control_external_wAddr_0) begin
          dataRegister_14 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'he == io_control_internal_wAddr_0) begin
              dataRegister_14 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'he == io_control_internal_wAddr_0) begin
            dataRegister_14 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_15 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'hf == io_control_external_wAddr_0) begin
          dataRegister_15 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'hf == io_control_internal_wAddr_0) begin
              dataRegister_15 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'hf == io_control_internal_wAddr_0) begin
            dataRegister_15 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_16 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h10 == io_control_external_wAddr_0) begin
          dataRegister_16 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h10 == io_control_internal_wAddr_0) begin
              dataRegister_16 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h10 == io_control_internal_wAddr_0) begin
            dataRegister_16 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_17 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h11 == io_control_external_wAddr_0) begin
          dataRegister_17 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h11 == io_control_internal_wAddr_0) begin
              dataRegister_17 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h11 == io_control_internal_wAddr_0) begin
            dataRegister_17 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_18 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h12 == io_control_external_wAddr_0) begin
          dataRegister_18 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h12 == io_control_internal_wAddr_0) begin
              dataRegister_18 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h12 == io_control_internal_wAddr_0) begin
            dataRegister_18 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_19 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h13 == io_control_external_wAddr_0) begin
          dataRegister_19 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h13 == io_control_internal_wAddr_0) begin
              dataRegister_19 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h13 == io_control_internal_wAddr_0) begin
            dataRegister_19 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_20 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h14 == io_control_external_wAddr_0) begin
          dataRegister_20 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h14 == io_control_internal_wAddr_0) begin
              dataRegister_20 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h14 == io_control_internal_wAddr_0) begin
            dataRegister_20 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_21 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h15 == io_control_external_wAddr_0) begin
          dataRegister_21 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h15 == io_control_internal_wAddr_0) begin
              dataRegister_21 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h15 == io_control_internal_wAddr_0) begin
            dataRegister_21 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_22 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h16 == io_control_external_wAddr_0) begin
          dataRegister_22 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h16 == io_control_internal_wAddr_0) begin
              dataRegister_22 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h16 == io_control_internal_wAddr_0) begin
            dataRegister_22 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_23 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h17 == io_control_external_wAddr_0) begin
          dataRegister_23 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h17 == io_control_internal_wAddr_0) begin
              dataRegister_23 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h17 == io_control_internal_wAddr_0) begin
            dataRegister_23 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_24 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h18 == io_control_external_wAddr_0) begin
          dataRegister_24 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h18 == io_control_internal_wAddr_0) begin
              dataRegister_24 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h18 == io_control_internal_wAddr_0) begin
            dataRegister_24 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_25 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h19 == io_control_external_wAddr_0) begin
          dataRegister_25 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h19 == io_control_internal_wAddr_0) begin
              dataRegister_25 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h19 == io_control_internal_wAddr_0) begin
            dataRegister_25 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_26 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h1a == io_control_external_wAddr_0) begin
          dataRegister_26 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h1a == io_control_internal_wAddr_0) begin
              dataRegister_26 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h1a == io_control_internal_wAddr_0) begin
            dataRegister_26 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_27 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h1b == io_control_external_wAddr_0) begin
          dataRegister_27 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h1b == io_control_internal_wAddr_0) begin
              dataRegister_27 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h1b == io_control_internal_wAddr_0) begin
            dataRegister_27 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_28 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h1c == io_control_external_wAddr_0) begin
          dataRegister_28 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h1c == io_control_internal_wAddr_0) begin
              dataRegister_28 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h1c == io_control_internal_wAddr_0) begin
            dataRegister_28 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_29 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h1d == io_control_external_wAddr_0) begin
          dataRegister_29 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h1d == io_control_internal_wAddr_0) begin
              dataRegister_29 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h1d == io_control_internal_wAddr_0) begin
            dataRegister_29 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_30 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h1e == io_control_external_wAddr_0) begin
          dataRegister_30 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h1e == io_control_internal_wAddr_0) begin
              dataRegister_30 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h1e == io_control_internal_wAddr_0) begin
            dataRegister_30 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      dataRegister_31 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        if (5'h1f == io_control_external_wAddr_0) begin
          dataRegister_31 <= io_wExternal_0;
        end else begin
          if (io_control_internal_wEnable_0) begin
            if (5'h1f == io_control_internal_wAddr_0) begin
              dataRegister_31 <= io_wInternal_0;
            end
          end
        end
      end else begin
        if (io_control_internal_wEnable_0) begin
          if (5'h1f == io_control_internal_wAddr_0) begin
            dataRegister_31 <= io_wInternal_0;
          end
        end
      end
    end
    if (reset) begin
      bpRegisterInt_0 <= 8'sh0;
    end else begin
      if (io_control_internal_wEnable_0) begin
        bpRegisterInt_0 <= io_wInternal_0;
      end
    end
    if (reset) begin
      bpRegisterExt_0 <= 8'sh0;
    end else begin
      if (io_control_external_wEnable_0) begin
        bpRegisterExt_0 <= io_wExternal_0;
      end
    end
  end
endmodule
